module Shift(A,B,ALUFun,S);
  input [31:0] A,B;
  input [5:0] ALUFun;//[1:0]
  output reg[31:0] S;
  
  wire [4:0] a;
  wire[31:0] b,c;
  reg [31:0] s0,s1,s2,s3;
  
  assign a=A[4:0];
  assign  b=0;
  assign  c=~b;

 
  
  always @(*) begin
    case(ALUFun[1:0])
      2'b00:begin
        s0=(a[0]==0)?B:{B[30:0],b[0]};
        s1=(a[1]==0)?s0:{s0[29:0],b[1:0]};
        s2=(a[2]==0)?s1:{s1[27:0],b[3:0]};
        s3=(a[3]==0)?s2:{s2[23:0],b[7:0]};
        S=(a[4]==0)?s3:{s3[15:0],b[15:0]};
      end
      2'b01:begin
        s0=(a[0]==0)?B:{b[31],B[31:1]};//1
        s1=(a[1]==0)?s0:{b[31:30],s0[31:2]};//2
        s2=(a[2]==0)?s1:{b[31:28],s1[31:4]};//4
        s3=(a[3]==0)?s2:{b[31:24],s2[31:8]};//8
        S=(a[4]==0)?s3:{b[31:16],s3[31:16]};//16
      end
      2'b11:begin
        case(B[31])
          1'b0:begin 
              s0=(a[0]==0)?B:{b[31],B[31:1]};//1
              s1=(a[1]==0)?s0:{b[31:30],s0[31:2]};//2
              s2=(a[2]==0)?s1:{b[31:28],s1[31:4]};//4
              s3=(a[3]==0)?s2:{b[31:24],s2[31:8]};//8
              S=(a[4]==0)?s3:{b[31:6],s3[31:16]};//16
              end
          1'b1:begin
              s0=(a[0]==0)?B:{c[31],B[31:1]};//1
              s1=(a[1]==0)?s0:{c[31:30],s0[31:2]};//2
              s2=(a[2]==0)?s1:{c[31:28],s1[31:4]};//4
              s3=(a[3]==0)?s2:{c[31:24],s2[31:8]};//8
              S=(a[4]==0)?s3:{c[31:16],s3[31:16]};//16
              end
            endcase
          end
    endcase
end
endmodule
  
  